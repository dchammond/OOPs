module cache
#(
)
(
);
endmodule : cache
